entity life_signs is
end;
